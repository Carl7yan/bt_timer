../../../common/8ut/tc/tc_1.sv