../../common/8ut/tb.sv