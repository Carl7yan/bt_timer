module tb;
  bit pclk;
  bit presetn;
  bit pclkg;

  initial begin
    forever
  end

cmsdk_apb_timer dut

endmodule