// ===================================================================
// Copyright (c) 2023 Carl Yan
// Owner      : carl.shengjie.yan@gmail.com
// Date       :
// Filename   :
// Abstract   :
//
// ===================================================================

// ===================================================================
// initial
initial begin
  #1_000_000  $finish;
end

// ===================================================================
// assertion
`ifdef SOC_ASSERT_ON

`endif
