// ===================================================================
// Copyright (c) 2023 Carl Yan
// Owner      : carl.shengjie.yan@gmail.com
// Date       :
// Filename   :
// Abstract   :
//
// ===================================================================

// ===================================================================
// initial
initial begin
  #2000  $finish;
end

// ===================================================================
// assertion
`ifdef SOC_ASSERT_ON

`endif
